module block_column (

);



endmodule