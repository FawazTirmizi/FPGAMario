module block_array (
    input logic Clk, Reset 
);

endmodule