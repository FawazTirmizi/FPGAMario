module FPGAMario_toplevel (

);

// big progresses lets gooooooo

endmodule